module balanced_less
(
   input [15:0] a, b, output q
);
   assign q = a < b; // TODO: check tree reported as balanced tree and not as ripple chain

endmodule
